grammar edu:umn:cs:melt:exts:ableC:wuffs;

exports edu:umn:cs:melt:exts:ableC:wuffs:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:wuffs:concretesyntax;
