grammar edu:umn:cs:melt:exts:ableC:asyncIO:concretesyntax;

terminal Spawn_t 'spawn' lexer classes {Keyword};
