grammar edu:umn:cs:melt:exts:ableC:asyncIO:concretesyntax;

terminal Spawn_t 'spawn' lexer classes {Keyword};
terminal Await_t 'await' lexer classes {Keyword};
