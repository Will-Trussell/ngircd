grammar edu:umn:cs:melt:exts:ableC:asyncIO;

exports edu:umn:cs:melt:exts:ableC:asyncIO:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:asyncIO:concretesyntax;
